module wzip

interface IWZipFile {
	path string
}
