module wzip

interface WZipFile {
	path string
}
